module video( );






endmodule
